-- 4-bit RGB values for VGA output

library ieee;
use ieee.std_logic_1164.all;

package stack_pkg is
    
end package stack_pkg;