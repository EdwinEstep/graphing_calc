entity alu is

end alu;